module top;
    initial begin

    end
endmodule : top
