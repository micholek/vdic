class env extends uvm_env;

    `uvm_component_utils(env)

    random_tester random_tester_h;
    driver driver_h;
    uvm_tlm_fifo#(alu_input_t) alu_input_f;

    coverage coverage_h;
    scoreboard scoreboard_h;
    alu_input_monitor alu_input_monitor_h;
    result_monitor result_monitor_h;

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction : new

    function void build_phase(uvm_phase phase);
        alu_input_f = new("alu_input_f", this);
        random_tester_h = random_tester::type_id::create("random_tester_h", this);
        driver_h = driver::type_id::create("drive_h", this);
        coverage_h = coverage::type_id::create ("coverage_h", this);
        scoreboard_h = scoreboard::type_id::create("scoreboard_h", this);
        alu_input_monitor_h = alu_input_monitor::type_id::create("alu_input_monitor_h", this);
        result_monitor_h = result_monitor::type_id::create("result_monitor_h", this);
    endfunction : build_phase

    function void connect_phase(uvm_phase phase);
        driver_h.alu_input_port.connect(alu_input_f.get_export);
        random_tester_h.alu_input_port.connect(alu_input_f.put_export);
        result_monitor_h.ap.connect(scoreboard_h.analysis_export);
        alu_input_monitor_h.ap.connect(scoreboard_h.alu_input_f.analysis_export);
        alu_input_monitor_h.ap.connect(coverage_h.analysis_export);
    endfunction : connect_phase

    function void end_of_elaboration_phase(uvm_phase phase);
        super.end_of_elaboration_phase(phase);
        $write("\033\[1;30m\033\[103m");
        $write("*** Created tester type: %s", random_tester_h.get_type_name());
        $write("\033\[0m\n");
    endfunction : end_of_elaboration_phase

endclass : env
